module uart_top()